magic
tech sky130B
magscale 1 2
timestamp 1719596937
<< error_s >>
rect 1070 600 1076 606
rect 1064 594 1070 600
rect 1064 540 1070 546
rect 1070 534 1076 540
rect 973 210 990 218
rect 1074 210 1120 218
rect 1204 210 1250 218
rect 1744 210 1790 218
rect 1874 210 1920 218
rect 2004 210 2050 218
rect 2544 210 2590 218
rect 2674 210 2720 218
rect 2804 210 2850 218
rect 3344 210 3390 218
rect 3474 210 3520 218
rect 3604 210 3650 218
rect 4144 210 4190 218
rect 4274 210 4320 218
rect 4404 210 4450 218
rect 4944 210 4990 218
rect 5074 210 5120 218
rect 5204 210 5237 218
rect 1001 182 1018 190
rect 1046 182 1148 190
rect 1176 182 1278 190
rect 1716 182 1818 190
rect 1846 182 1948 190
rect 1976 182 2078 190
rect 2516 182 2618 190
rect 2646 182 2748 190
rect 2776 182 2878 190
rect 3316 182 3418 190
rect 3446 182 3548 190
rect 3576 182 3678 190
rect 4116 182 4218 190
rect 4246 182 4348 190
rect 4376 182 4478 190
rect 4916 182 5018 190
rect 5046 182 5148 190
rect 5176 182 5209 190
<< locali >>
rect 860 400 960 740
rect 1240 400 1340 740
rect 1660 400 1760 740
rect 2040 400 2140 740
rect 2460 400 2560 740
rect 2840 400 2940 740
rect 3260 400 3360 740
rect 3640 400 3740 740
rect 4060 400 4160 740
rect 4440 400 4540 740
rect 4860 400 4960 740
rect 5240 400 5340 740
rect 880 0 1320 40
rect 1680 0 2120 40
rect 2480 0 2920 40
rect 3280 0 3720 40
rect 4080 0 4520 40
rect 4880 0 5320 40
rect 800 -100 5400 0
<< metal1 >>
rect 1001 960 5209 1019
rect 1870 600 1930 606
rect 1060 540 1070 600
rect 1130 540 1140 600
rect 1870 534 1930 540
rect 2670 600 2730 606
rect 2670 534 2730 540
rect 4270 600 4330 606
rect 4270 534 4330 540
rect 5070 600 5130 606
rect 5070 534 5130 540
rect 1001 131 5209 190
<< via1 >>
rect 1070 540 1130 600
rect 1870 540 1930 600
rect 2670 540 2730 600
rect 4270 540 4330 600
rect 5070 540 5130 600
<< metal2 >>
rect 1130 540 1870 600
rect 1930 540 2670 600
rect 2730 540 4270 600
rect 4330 540 5070 600
rect 5130 540 5136 600
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_0
timestamp 1719596467
transform 1 0 5097 0 1 570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_1
timestamp 1719596467
transform 1 0 1097 0 1 570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_2
timestamp 1719596467
transform 1 0 1897 0 1 570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_3
timestamp 1719596467
transform 1 0 2697 0 1 570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_4
timestamp 1719596467
transform 1 0 3497 0 1 570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_5
timestamp 1719596467
transform 1 0 4297 0 1 570
box -297 -570 297 570
<< end >>
